module platform2(
    input wire p2_on,			// signal from colour sensor module to initiate platform2 module
    input wire clk,     		// 50 MHz
    input wire [5:0] colour, 		// colour data input from colour sensor
    output reg [3:0] GPIO_1,		// output to the physical motor turning the platform (1st motor)
    output reg motor_on			// output to "motor" module (that controls the 2nd motor)
);
	 
motor motor_(.motor_on(motor_on));
	
// Stores the input signal of p2_on(1) and allows it to changed back to 0
reg p2_on_internal;
	
// Controls speed of motor
reg [31:0] count = 390_624;  

// Controls timing of motor
reg [31:0] cntr = 0;

// Controls the number of clock cycles the motor runs for
// 1 full rotation = 50 mill, given a 50MHs clock
reg [31:0] timer = 50_000_000;

// Clockwise locations
reg [31:0] red_timer = (50_000_000 * 0.125); // Red location    = 45/360
reg [31:0] bro_timer = (50_000_000 * 0.250); // Brown location  = 90/360
reg [31:0] yel_timer = (50_000_000 * 0.375); // Yellow location = 135/360
reg [31:0] ora_timer = (50_000_000 * 0.500); // Orange location = 180/360

// Counter clockwise locations
reg [31:0] blu_timer = (50_000_000 * 0.250); // Blue location   = 90/360
reg [31:0] gre_timer = (50_000_000 * 0.375); // Green location  = 135/360

always @(posedge clk) begin
    p2_on_internal <= p2_on; 		// Store p2_on signal

    if (p2_on_internal == 1) begin 	// Check if p2 module ready to begin
    
    p2_on_internal <= 0; 		// Then change back to 0

    // RED Begin
    if (colour == 000001) begin
    if (red_timer > 0) begin
        if (cntr < count*1/4) begin
            GPIO_1 <= 4'b1000;
        end else if (cntr < count*2/4) begin
            GPIO_1 <= 4'b0100;
        end else if (cntr < count*3/4) begin
            GPIO_1 <= 4'b0010;
        end else if (cntr < count*4/4) begin
            GPIO_1 <= 4'b0001;
        red_timer <= red_timer - 1; // Countdown to zero
        end
        cntr <= cntr + 1;
        if (cntr >= count) begin
            cntr <= 0;
        end  
        end else begin
        GPIO_1 <= 4'b0000; 	 // M&M is above it's respective colour bin - stop motor
        motor_on <= 1;		 // Call Motor module to open latch and let M&M fall into bin
        end
    end // RED end

    // BROWN Begin
    else if (colour == 000010) begin
    if (bro_timer > 0) begin
        if (cntr < count*1/4) begin
            GPIO_1 <= 4'b1000;
        end else if (cntr < count*2/4) begin
            GPIO_1 <= 4'b0100;
        end else if (cntr < count*3/4) begin
            GPIO_1 <= 4'b0010;
        end else if (cntr < count*4/4) begin
            GPIO_1 <= 4'b0001;
        bro_timer <= bro_timer - 1; // Countdown to zero
        end
        cntr <= cntr + 1;
        if (cntr >= count) begin
            cntr <= 0;
        end  
        end else begin
        GPIO_1 <= 4'b0000; 	 // M&M is above it's respective colour bin - stop motor
        motor_on <= 1;		 // Call Motor module to open latch and let M&M fall into bin
        end
    end // Brown end

    // YELLOW Begin
    else if (colour == 000100) begin
    if (yel_timer > 0) begin
        if (cntr < count*1/4) begin
            GPIO_1 <= 4'b1000;
        end else if (cntr < count*2/4) begin
            GPIO_1 <= 4'b0100;
        end else if (cntr < count*3/4) begin
            GPIO_1 <= 4'b0010;
        end else if (cntr < count*4/4) begin
            GPIO_1 <= 4'b0001;
        yel_timer <= yel_timer - 1; // Countdown to zero
        end
        cntr <= cntr + 1;
        if (cntr >= count) begin
            cntr <= 0;
        end  
        end else begin
        GPIO_1 <= 4'b0000; 	 // M&M is above it's respective colour bin - stop motor
        motor_on <= 1;		 // Call Motor module to open latch and let M&M fall into bin
        end
    end // Yellow end

    // ORANGE Begin
    else if (colour == 001000) begin
    if (ora_timer > 0) begin
        if (cntr < count*1/4) begin
            GPIO_1 <= 4'b1000;
        end else if (cntr < count*2/4) begin
            GPIO_1 <= 4'b0100;
        end else if (cntr < count*3/4) begin
            GPIO_1 <= 4'b0010;
        end else if (cntr < count*4/4) begin
            GPIO_1 <= 4'b0001;
        ora_timer <= ora_timer - 1; // Countdown to zero
        end
        cntr <= cntr + 1;
        if (cntr >= count) begin
            cntr <= 0;
        end  
        end else begin
        GPIO_1 <= 4'b0000; 	 // M&M is above it's respective colour bin - stop motor
        motor_on <= 1;		 // Call Motor module to open latch and let M&M fall into bin
        end
    end // Orange end

    // BLUE Begin
    else if (colour == 010000) begin
    if (blu_timer > 0) begin
        if (cntr < count*1/4) begin
            GPIO_1 <= 4'b0001;
        end else if (cntr < count*2/4) begin
            GPIO_1 <= 4'b0010;
        end else if (cntr < count*3/4) begin
            GPIO_1 <= 4'b0100;
        end else if (cntr < count*4/4) begin
            GPIO_1 <= 4'b1000;
        blu_timer <= blu_timer - 1; // Countdown to zero
        end
        cntr <= cntr + 1;
        if (cntr >= count) begin
            cntr <= 0;
        end  
        end else begin
        GPIO_1 <= 4'b0000; 	 // M&M is above it's respective colour bin - stop motor
        motor_on <= 1;		 // Call Motor module to open latch and let M&M fall into bin
        end
    end // Blue end

    // GREEN Begin
    else if (colour == 100000) begin
    if (gre_timer > 0) begin
        if (cntr < count*1/4) begin
            GPIO_1 <= 4'b0001;
        end else if (cntr < count*2/4) begin
            GPIO_1 <= 4'b0010;
        end else if (cntr < count*3/4) begin
            GPIO_1 <= 4'b0100;
        end else if (cntr < count*4/4) begin
            GPIO_1 <= 4'b1000;
        gre_timer <= gre_timer - 1; // Countdown to zero
        end
        cntr <= cntr + 1;
        if (cntr >= count) begin
            cntr <= 0;
        end  
        end else begin
        GPIO_1 <= 4'b0000; 	 // M&M is above it's respective colour bin - stop motor
        motor_on <= 1;		 // Call Motor module to open latch and let M&M fall into bin
        end
    end // Green end
  end // motor_on end
end // clk end
endmodule
